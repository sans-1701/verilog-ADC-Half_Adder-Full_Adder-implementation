module 4_Bit_Op(
    input wire [3:0] A , B ; 
    input wire T ; 
    output wire [3:0] S;
    output wire Cout;
);